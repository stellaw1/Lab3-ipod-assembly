
`default_nettype none
 `define USE_PACOBLAZE
module 
picoblaze_template
#(
parameter clk_freq_in_hz = 25000000
) (
  output reg[7:0] led,
  output reg led0,
  input clk, interrupt_event, 
  input [7:0] input_data,
  output wire [23:0] sseg
);

  
//--
//------------------------------------------------------------------------------------
//--
//-- Signals used to connect KCPSM3 to program ROM and I/O logic
//--

wire[9:0]  address;
wire[17:0]  instruction;
wire[7:0]  port_id;
wire[7:0]  out_port;
reg[7:0]  in_port;
wire  write_strobe;
wire  read_strobe;
reg  interrupt;
wire  interrupt_ack;
wire  kcpsm3_reset;


//-- Signals for LCD operation
//--
//--

reg        lcd_rw_control;
reg[7:0]   lcd_output_data;
pacoblaze3 led_8seg_kcpsm
(
                  .address(address),
               .instruction(instruction),
                   .port_id(port_id),
              .write_strobe(write_strobe),
                  .out_port(out_port),
               .read_strobe(read_strobe),
                   .in_port(in_port),
                 .interrupt(interrupt),
             .interrupt_ack(interrupt_ack),
                     .reset(kcpsm3_reset),
                       .clk(clk));

wire [19:0] raw_instruction;

pacoblaze_instruction_memory 
pacoblaze_instruction_memory_inst(
  .addr(address),
  .outdata(raw_instruction)
);

always @ (posedge clk)
begin
  instruction <= raw_instruction[17:0];
end

assign kcpsm3_reset = 0;                       
  
//  ----------------------------------------------------------------------------------------------------------------------------------
//  -- Interrupt 
//  ----------------------------------------------------------------------------------------------------------------------------------
//  --
//  --
//  -- Interrupt is used to provide a 1 second time reference.
//  --
//  --
//  -- A simple binary counter is used to divide the 50MHz system clock and provide interrupt pulses.
//  --


// Note that because we are using clock enable we DO NOT need to synchronize with clk

always @ (posedge clk or posedge interrupt_ack)  //FF with clock "clk" and reset "interrupt_ack"
begin
  if (interrupt_ack) //if we get reset, reset interrupt in order to wait for next clock.
    interrupt <= 0;
  else
begin 
  if (interrupt_event)   //clock enable
    interrupt <= 1;
  else
    interrupt <= interrupt;
  end
end

//  --
//  ----------------------------------------------------------------------------------------------------------------------------------
//  -- KCPSM3 input ports 
//  ----------------------------------------------------------------------------------------------------------------------------------
//  --
//  --
//  -- The inputs connect via a pipelined multiplexer
//  --

always @ (posedge clk)
begin
  case (port_id[7:0])
    8'h0:    in_port <= input_data;
    default: in_port <= 8'bx;
  endcase
end
   
//
//  --
//  ----------------------------------------------------------------------------------------------------------------------------------
//  -- KCPSM3 output ports 
//  ----------------------------------------------------------------------------------------------------------------------------------
//  --
//  -- adding the output registers to the processor
//  --
//   
always @ (posedge clk)
begin

  //port 80 hex 
  if (write_strobe & port_id[7])  //clock enable 
    led <= out_port;

  //port 40 hex 
  if (write_strobe & port_id[6])  //clock enable 
    sseg[7:0] <= out_port;
      
  //port 20 hex 
  if (write_strobe & port_id[5])  //clock enable 
    sseg[15:8] <= out_port;
      
  //port 10 hex 			
  if (write_strobe & port_id[4])  //clock enable 
    sseg[23:16] <= out_port;
  
  //port 8 hex 			
  if (write_strobe & port_id[3])  //clock enable 
    led0 <= out_port;
          
end

endmodule
